

module fwuart(
);

endmodule

